// Lookup table for function log((1+e^(-|x|)) / (1-e^(-|x|)) )
// X: 6 bits, 2 integer: 4 fractional, thus can be sampled at 0.0625
// Y: 4 bits, 2 integer: 2 fractional, thus can be quantized at 0.25

module LUT (
  input [6-1 : 0] X,
  output reg [4-1 : 0] Y
);

always@ (X) begin
  case (X)
    6'b000000: Y = 4'b1111;  // f(0.0)   = 3.75 ~ 3.75
    6'b000001: Y = 4'b1000;  // f(0.25)  = 2.0846309693248757 ~ 2.0
    6'b000010: Y = 4'b0110;  // f(0.5)   = 1.4068291137472952 ~ 1.5
    6'b000011: Y = 4'b0100;  // f(0.75)  = 1.0262244711552542 ~ 1.0
    6'b000100: Y = 4'b0011;  // f(1.0)   = 0.7719368329053048 ~ 0.75
    6'b000101: Y = 4'b0010;  // f(1.25)  = 0.589508646432784 ~ 0.5
    6'b000110: Y = 4'b0010;  // f(1.5)   = 0.4538957369082066 ~ 0.5
    6'b000111: Y = 4'b0001;  // f(1.75)  = 0.3511110171316341 ~ 0.25
    6'b001000: Y = 4'b0001;  // f(2.0)   = 0.2723414689118317 ~ 0.25
    6'b001001: Y = 4'b0001;  // f(2.25)  = 0.21158428010179142 ~ 0.25
    6'b001010: Y = 4'b0001;  // f(2.5)   = 0.1645402180345878 ~ 0.25
    6'b001011: Y = 4'b0001;  // f(2.75)  = 0.1280303231172332 ~ 0.25
    6'b001100: Y = 4'b0000;  // f(3.0)   = 0.09965653251644369 ~ 0.0
    6'b001101: Y = 4'b0000;  // f(3.25)  = 0.077587313867282 ~ 0.0
    6'b001110: Y = 4'b0000;  // f(3.5)   = 0.06041313452808037 ~ 0.0
    6'b001111: Y = 4'b0000;  // f(3.75)  = 0.0470441661225781 ~ 0.0
    6'b010000: Y = 4'b0000;  // f(4.0)   = 0.03663537474369636 ~ 0.0
    6'b010001: Y = 4'b0000;  // f(4.25)  = 0.028530402934517397 ~ 0.0
    6'b010010: Y = 4'b0000;  // f(4.5)   = 0.02221890711689061 ~ 0.0
    6'b010011: Y = 4'b0000;  // f(4.75)  = 0.017303822155776718 ~ 0.0
    6'b010100: Y = 4'b0000;  // f(5.0)   = 0.013476097938606508 ~ 0.0
    6'b010101: Y = 4'b0000;  // f(5.25)  = 0.010495133131970643 ~ 0.0
    6'b010110: Y = 4'b0000;  // f(5.5)   = 0.008173588381406572 ~ 0.0
    6'b010111: Y = 4'b0000;  // f(5.75)  = 0.006365583087728265 ~ 0.0
    6'b011000: Y = 4'b0000;  // f(6.0)   = 0.0049575145066898104 ~ 0.0
    6'b011001: Y = 4'b0000;  // f(6.25)  = 0.003860913068554783 ~ 0.0
    6'b011010: Y = 4'b0000;  // f(6.5)   = 0.003006880651470039 ~ 0.0
    6'b011011: Y = 4'b0000;  // f(6.75)  = 0.002341760311735284 ~ 0.0
    6'b011100: Y = 4'b0000;  // f(7.0)   = 0.001823764436613251 ~ 0.0
    6'b011101: Y = 4'b0000;  // f(7.25)  = 0.0014203490164682224 ~ 0.0
    6'b011110: Y = 4'b0000;  // f(7.5)   = 0.0011061688530888379 ~ 0.0
    6'b011111: Y = 4'b0000;  // f(7.75)  = 0.0008614851344310268 ~ 0.0
    6'b100000: Y = 4'b0000;  // f(8.0)   = 0.000670925280972407 ~ 0.0
    6'b100001: Y = 4'b0000;  // f(8.25)  = 0.0005225171264915748 ~ 0.0
    6'b100010: Y = 4'b0000;  // f(8.5)   = 0.00040693674363700874 ~ 0.0
    6'b100011: Y = 4'b0000;  // f(8.75)  = 0.00031692265288412293 ~ 0.0
    6'b100100: Y = 4'b0000;  // f(9.0)   = 0.0002468196094264098 ~ 0.0
    6'b100101: Y = 4'b0000;  // f(9.25)  = 0.00019222330471475586 ~ 0.0
    6'b100110: Y = 4'b0000;  // f(9.5)   = 0.00014970366005496292 ~ 0.0
    6'b100111: Y = 4'b0000;  // f(9.75)  = 0.00011658932759383428 ~ 0.0
    6'b101000: Y = 4'b0000;  // f(10.0)  = 9.079985958730571e-05 ~ 0.0
    6'b101001: Y = 4'b0000;  // f(10.25) = 7.071500173041337e-05 ~ 0.0
    6'b101010: Y = 4'b0000;  // f(10.5)  = 5.507289871350473e-05 ~ 0.0
    6'b101011: Y = 4'b0000;  // f(10.75) = 4.289081663965259e-05 ~ 0.0
    6'b101100: Y = 4'b0000;  // f(11.0)  = 3.3403401583538476e-05 ~ 0.0
    6'b101101: Y = 4'b0000;  // f(11.25) = 2.60145953096234e-05 ~ 0.0
    6'b101110: Y = 4'b0000;  // f(11.5)  = 2.0260187197876252e-05 ~ 0.0
    6'b101111: Y = 4'b0000;  // f(11.75) = 1.577864965483916e-05 ~ 0.0
    6'b110000: Y = 4'b0000;  // f(12.0)  = 1.2288424706844796e-05 ~ 0.0
    6'b110001: Y = 4'b0000;  // f(12.25) = 9.570234784286784e-06 ~ 0.0
    6'b110010: Y = 4'b0000;  // f(12.5)  = 7.453306344154328e-06 ~ 0.0
    6'b110011: Y = 4'b0000;  // f(12.75) = 5.804640817349936e-06 ~ 0.0
    6'b110100: Y = 4'b0000;  // f(13.0)  = 4.520658814032911e-06 ~ 0.0
    6'b110101: Y = 4'b0000;  // f(13.25) = 3.5206926241672784e-06 ~ 0.0
    6'b110110: Y = 4'b0000;  // f(13.5)  = 2.74191817288693e-06 ~ 0.0
    6'b110111: Y = 4'b0000;  // f(13.75) = 2.1354080201560868e-06 ~ 0.0
    6'b111000: Y = 4'b0000;  // f(14.0)  = 1.6630574382189508e-06 ~ 0.0
    6'b111001: Y = 4'b0000;  // f(14.25) = 1.2951904352494061e-06 ~ 0.0
    6'b111010: Y = 4'b0000;  // f(14.5)  = 1.008695325015218e-06 ~ 0.0
    6'b111011: Y = 4'b0000;  // f(14.75) = 7.85572709185188e-07 ~ 0.0
    6'b111100: Y = 4'b0000;  // f(15.0)  = 6.11804640979781e-07 ~ 0.0
    6'b111101: Y = 4'b0000;  // f(15.25) = 4.7647393359265615e-07 ~ 0.0
    6'b111110: Y = 4'b0000;  // f(15.5)  = 3.710782725383919e-07 ~ 0.0
    6'b111111: Y = 4'b0000;  // f(15.75) = 2.889960492985625e-07 ~ 0.0
    default:   Y = 0;
  endcase

end

endmodule
